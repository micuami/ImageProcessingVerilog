module test_image1;

tester tester();

endmodule

